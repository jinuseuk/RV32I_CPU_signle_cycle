`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);

    logic [31:0] rom[0:2**8-1];

    initial begin
     
        rom[0] = 32'b0000000_00001_00010_000_00100_0110011;  // add x4, x2, x1 (x4 = x2 + x1)
        rom[1] = 32'b0100000_00001_00010_000_00101_0110011;  // sub x5, x2, x1 (x5 = x2 - x1)
        rom[2] = 32'b0000000_00000_00011_111_00110_0110011;  // and x6, x3, x0 (x6 = x3 & x0)
        rom[3] = 32'b0000000_00000_00011_110_00111_0110011;  // or  x7, x3, x0 (x7 = x3 | x0)
        

        rom[4] = 32'b0000000_00010_00011_100_01000_0110011;  // xor x8, x3, x2
        rom[5] = 32'b0000000_00001_00100_001_01001_0110011;  // sll x9, x4, x1
        rom[6] = 32'b0000000_00010_00011_010_01010_0110011;  // slt x10, x3, x2 (부호있는 비교)
        rom[7] = 32'b0000000_00011_00010_011_01011_0110011;  // sltu x11, x2, x3 (부호없는 비교)
        rom[8] = 32'b0000000_00001_00100_101_01100_0110011;  // srl x12, x4, x1
        rom[9] = 32'b0100000_00001_00100_101_01101_0110011;  // sra x13, x4, x1


   
        rom[10] = 32'b000000000001_00001_000_01001_0010011;  // addi x9, x1, 1 (원래 rom[4])
        rom[11] = 32'b000000000100_00010_111_01010_0010011;  // andi x10, x2, 4 (원래 rom[5])
        rom[12] = 32'b000000000011_00001_001_01011_0010011;  // slli x11, x1, 3 (원래 rom[6])
        rom[13] = 32'b000000001001_00001_001_01100_0010011;  // slli x12, x1, 9 (원래 rom[7])
        rom[14] = 32'b000000011110_00001_001_01101_0010011;  // slli x13, x1, 30 (원래 rom[8])

     
        rom[15] = 32'b111111111100_00010_100_01110_0010011;  // xori x14, x2, -4 (음수 즉치값 테스트)
        rom[16] = 32'b000000000111_00011_110_01111_0010011;  // ori x15, x3, 7
        rom[17] = 32'b000000000101_00100_010_10000_0010011;  // slti x16, x4, 5
        rom[18] = 32'b0000000_00000_00101_101_10001_0010011;  // srli x17, x5, 0 (rs1=x5, shamt=0, Funct7=0000000)
        rom[19] = 32'b0100000_00100_00101_101_10010_0010011;  // srai x18, x5, 4 (rs1=x5, shamt=4, Funct7=0100000)


        // [31:20] Imm _ [19:15] rs1 _ [14:12] Funct3 _ [11:7] rd _ [6:0] Opcode
        rom[20] = 32'b000000000100_00000_000_01110_0000011;  // lb x14, 4(x0) (원래 rom[15])
        rom[21] = 32'b000000001000_00000_001_01111_0000011;  // lh x15, 8(x0) (원래 rom[16])
        rom[22] = 32'b000000001100_00000_010_10000_0000011;  // lw x16, 12(x0) (원래 rom[17])

        rom[23] = 32'b000000010000_00000_100_10001_0000011;  // lbu x17, 16(x0) (Unsigned Byte Load)
        rom[24] = 32'b000000010100_00000_101_10010_0000011;  // lhu x18, 20(x0) (Unsigned Halfword Load)
        

 
        // [31:25] Imm[11:5] _ [24:20] rs2 _ [19:15] rs1 _ [14:12] Funct3 _ [11:7] Imm[4:0] _ [6:0] Opcode
        rom[25] = 32'b0000000_01011_00000_000_00100_0100011;  // sb x11, 4(x0) (원래 rom[12])
        rom[26] = 32'b0000000_01100_00000_001_01000_0100011;  // sh x12, 8(x0) (원래 rom[13])
        rom[27] = 32'b0000000_01101_00000_010_01100_0100011;  // sw x13, 12(x0) (원래 rom[14])
        
  
       
        // [31] Imm[12] _ [30:25] Imm[10:5] _ [24:20] rs2 _ [19:15] rs1 _ [14:12] Funct3 _ [11:8] Imm[4:1] _ [7] Imm[11] _ [6:0] Opcode
        rom[28] = 32'b0000000_00010_00010_000_01100_1100011;  // beq x2, x2, 12 (Branch to PC+12, 원래 rom[9])
        

        rom[29] = 32'b0000000_00010_00011_001_01000_1100011;  // bne x3, x2, 8 (Branch to PC+8)
        rom[30] = 32'b0000000_00010_00011_100_11000_1100011;  // blt x3, x2, 24 (Branch if x3 < x2)
        rom[31] = 32'b0000000_00011_00010_101_10100_1100011;  // bge x2, x3, 20 (Branch if x2 >= x3)
        rom[32] = 32'b0000000_00010_00011_110_10000_1100011;  // bltu x3, x2, 16 (Unsigned)
        rom[33] = 32'b0000000_00011_00010_111_10010_1100011;  // bgeu x2, x3, 18 (Unsigned)



        rom[34] = 32'b00010000000000000000_10001_0110111;  // lui x17, 0x100000 (원래 rom[18])
        

        rom[35] = 32'b00010000000000000000_10010_0010111;  // auipc x18, 0x100000 (PC + 0x100000 << 12)
        

        // [31] Imm[20] _ [30:21] Imm[10:1] _ [20] Imm[11] _ [19:12] Imm[19:12] _ [11:7] rd _ [6:0] Opcode
        rom[36] = 32'b00000001000000000000_00011_1101111;  // jal x3, 16 (Jump to PC+16, 원래 rom[17]의 LW와 충돌 방지 위해 이동)



        // [31:20] Imm _ [19:15] rs1 _ [14:12] Funct3 _ [11:7] rd _ [6:0] Opcode
        rom[37] = 32'b000000011100_00100_000_00100_1100111;  // jalr x4, 28(x4) (원래 rom[21])


        rom[38] = 32'b000000000000_00000_000_00000_0010011;  // addi x0, x0, 0
        rom[39] = 32'hFFFFFFFF;                               // Fill with FFFF (Stop/Halt Signal for Testbench)

    end


    assign data = rom[addr[31:2]];
endmodule
